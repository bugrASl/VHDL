library	IEEE;
use	IEEE.STD_LOGIC_1164.all;

package	parity_pkg	is
	type	PARITY_TYPE	is	(EVEN,ODD);
end	package;
